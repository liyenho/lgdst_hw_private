// altera_asmi.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module altera_asmi (
		input  wire [31:0] addr,       //       addr.addr
		output wire        busy,       //       busy.busy
		input  wire        clkin,      //      clkin.clk
		output wire        data_valid, // data_valid.data_valid
		output wire [7:0]  dataout,    //    dataout.dataout
		input  wire        en4b_addr,  //  en4b_addr.en4b_addr
		input  wire        rden,       //       rden.rden
		input  wire        read,       //       read.read
		input  wire        reset,      //      reset.reset
		input  wire        wren        //       wren.wren
	);

	altera_asmi_asmi_parallel_0 asmi_parallel_0 (
		.clkin      (clkin),      //      clkin.clk
		.read       (read),       //       read.read
		.rden       (rden),       //       rden.rden
		.addr       (addr),       //       addr.addr
		.wren       (wren),       //       wren.wren
		.en4b_addr  (en4b_addr),  //  en4b_addr.en4b_addr
		.reset      (reset),      //      reset.reset
		.dataout    (dataout),    //    dataout.dataout
		.busy       (busy),       //       busy.busy
		.data_valid (data_valid)  // data_valid.data_valid
	);

endmodule
