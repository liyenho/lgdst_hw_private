// system_bd.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module system_bd (
		input  wire         axi_ad9361_device_clock_clk,           //      axi_ad9361_device_clock.clk
		input  wire         axi_ad9361_device_if_rx_clk_in_p,      //         axi_ad9361_device_if.rx_clk_in_p
		input  wire         axi_ad9361_device_if_rx_clk_in_n,      //                             .rx_clk_in_n
		input  wire         axi_ad9361_device_if_rx_frame_in_p,    //                             .rx_frame_in_p
		input  wire         axi_ad9361_device_if_rx_frame_in_n,    //                             .rx_frame_in_n
		input  wire [5:0]   axi_ad9361_device_if_rx_data_in_p,     //                             .rx_data_in_p
		input  wire [5:0]   axi_ad9361_device_if_rx_data_in_n,     //                             .rx_data_in_n
		output wire         axi_ad9361_device_if_tx_clk_out_p,     //                             .tx_clk_out_p
		output wire         axi_ad9361_device_if_tx_clk_out_n,     //                             .tx_clk_out_n
		output wire         axi_ad9361_device_if_tx_frame_out_p,   //                             .tx_frame_out_p
		output wire         axi_ad9361_device_if_tx_frame_out_n,   //                             .tx_frame_out_n
		output wire [5:0]   axi_ad9361_device_if_tx_data_out_p,    //                             .tx_data_out_p
		output wire [5:0]   axi_ad9361_device_if_tx_data_out_n,    //                             .tx_data_out_n
		output wire         axi_ad9361_dma_if_adc_enable_i0,       //            axi_ad9361_dma_if.adc_enable_i0
		output wire         axi_ad9361_dma_if_adc_valid_i0,        //                             .adc_valid_i0
		output wire [15:0]  axi_ad9361_dma_if_adc_data_i0,         //                             .adc_data_i0
		output wire         axi_ad9361_dma_if_adc_enable_q0,       //                             .adc_enable_q0
		output wire         axi_ad9361_dma_if_adc_valid_q0,        //                             .adc_valid_q0
		output wire [15:0]  axi_ad9361_dma_if_adc_data_q0,         //                             .adc_data_q0
		output wire         axi_ad9361_dma_if_adc_enable_i1,       //                             .adc_enable_i1
		output wire         axi_ad9361_dma_if_adc_valid_i1,        //                             .adc_valid_i1
		output wire [15:0]  axi_ad9361_dma_if_adc_data_i1,         //                             .adc_data_i1
		output wire         axi_ad9361_dma_if_adc_enable_q1,       //                             .adc_enable_q1
		output wire         axi_ad9361_dma_if_adc_valid_q1,        //                             .adc_valid_q1
		output wire [15:0]  axi_ad9361_dma_if_adc_data_q1,         //                             .adc_data_q1
		input  wire         axi_ad9361_dma_if_adc_dovf,            //                             .adc_dovf
		input  wire         axi_ad9361_dma_if_adc_dunf,            //                             .adc_dunf
		output wire         axi_ad9361_dma_if_dac_enable_i0,       //                             .dac_enable_i0
		output wire         axi_ad9361_dma_if_dac_valid_i0,        //                             .dac_valid_i0
		input  wire [15:0]  axi_ad9361_dma_if_dac_data_i0,         //                             .dac_data_i0
		output wire         axi_ad9361_dma_if_dac_enable_q0,       //                             .dac_enable_q0
		output wire         axi_ad9361_dma_if_dac_valid_q0,        //                             .dac_valid_q0
		input  wire [15:0]  axi_ad9361_dma_if_dac_data_q0,         //                             .dac_data_q0
		output wire         axi_ad9361_dma_if_dac_enable_i1,       //                             .dac_enable_i1
		output wire         axi_ad9361_dma_if_dac_valid_i1,        //                             .dac_valid_i1
		input  wire [15:0]  axi_ad9361_dma_if_dac_data_i1,         //                             .dac_data_i1
		output wire         axi_ad9361_dma_if_dac_enable_q1,       //                             .dac_enable_q1
		output wire         axi_ad9361_dma_if_dac_valid_q1,        //                             .dac_valid_q1
		input  wire [15:0]  axi_ad9361_dma_if_dac_data_q1,         //                             .dac_data_q1
		input  wire         axi_ad9361_dma_if_dac_dovf,            //                             .dac_dovf
		input  wire         axi_ad9361_dma_if_dac_dunf,            //                             .dac_dunf
		output wire         axi_ad9361_master_if_l_clk,            //         axi_ad9361_master_if.l_clk
		input  wire         axi_ad9361_master_if_dac_sync_in,      //                             .dac_sync_in
		output wire         axi_ad9361_master_if_dac_sync_out,     //                             .dac_sync_out
		input  wire         axi_ad9361_user_if_usr_tx_data_sel,    //           axi_ad9361_user_if.usr_tx_data_sel
		input  wire [5:0]   axi_ad9361_user_if_usr_tx_data_i,    //                             .usr_tx_p_data_p
		input  wire [5:0]   axi_ad9361_user_if_usr_tx_data_q,    //                             .usr_tx_p_data_n
		input  wire         axi_ad9361_user_if_usr_tx_frame,     //                             .usr_tx_p_frame
		input  wire         clk_clk,                               //                          clk.clk
		output wire [4:0]   gpio_external_connection_export,       //     gpio_external_connection.export
		output wire         reg_map_usr_rd_word_en,                //                      reg_map.usr_rd_word_en
		output wire [7:0]   reg_map_usr_rd_word_addr,              //                             .usr_rd_word_addr
		input  wire [31:0]  reg_map_usr_rd_word_data,              //                             .usr_rd_word_data
		output wire         reg_map_usr_wr_word_en,                //                             .usr_wr_word_en
		output wire [3:0]   reg_map_usr_wr_byte_indx,              //                             .usr_wr_byte_indx
		output wire [7:0]   reg_map_usr_wr_word_addr,              //                             .usr_wr_word_addr
		output wire [31:0]  reg_map_usr_wr_word_data,              //                             .usr_wr_word_data
		output wire [255:0] reg_map_test_out,                      //                             .test_out
		input  wire         reset_reset_n,                         //                        reset.reset_n
		input  wire         spi_ad9361_external_MISO,              //          spi_ad9361_external.MISO
		output wire         spi_ad9361_external_MOSI,              //                             .MOSI
		output wire         spi_ad9361_external_SCLK,              //                             .SCLK
		output wire         spi_ad9361_external_SS_n,              //                             .SS_n
		input  wire [31:0]  sys_gpio_external_connection_in_port,  // sys_gpio_external_connection.in_port
		output wire [31:0]  sys_gpio_external_connection_out_port  //                             .out_port
	);

   pll_for_lvds i_pll_lvds(
    .refclk(axi_ad9361_device_if_rx_clk_in_p), 
    .rst(!reset_reset_n), 

    .outclk_0(axi_ad9361_device_if_tx_clk_out_p), 
    .outclk_1(axi_ad9361_device_if_tx_clk_out_n),
    .outclk_2(axi_ad9361_master_if_l_clk)
   );

endmodule
