// remote_update.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module remote_update (
		output wire [31:0] asmi_addr,       //       asmi_addr.asmi_addr
		input  wire        asmi_busy,       //       asmi_busy.asmi_busy
		input  wire        asmi_data_valid, // asmi_data_valid.asmi_data_valid
		input  wire [7:0]  asmi_dataout,    //    asmi_dataout.asmi_dataout
		output wire        asmi_rden,       //       asmi_rden.asmi_rden
		output wire        asmi_read,       //       asmi_read.asmi_read
		output wire        busy,            //            busy.busy
		input  wire        clock,           //           clock.clk
		input  wire [31:0] data_in,         //         data_in.data_in
		output wire [31:0] data_out,        //        data_out.data_out
		input  wire [2:0]  param,           //           param.param
		output wire        pof_error,       //       pof_error.pof_error
		input  wire        read_param,      //      read_param.read_param
		input  wire        reconfig,        //        reconfig.reconfig
		input  wire        reset,           //           reset.reset
		input  wire        reset_timer,     //     reset_timer.reset_timer
		input  wire        write_param      //     write_param.write_param
	);

	remote_update_remote_update_0 remote_update_0 (
		.busy            (busy),            //            busy.busy
		.data_out        (data_out),        //        data_out.data_out
		.param           (param),           //           param.param
		.read_param      (read_param),      //      read_param.read_param
		.reconfig        (reconfig),        //        reconfig.reconfig
		.reset_timer     (reset_timer),     //     reset_timer.reset_timer
		.write_param     (write_param),     //     write_param.write_param
		.data_in         (data_in),         //         data_in.data_in
		.clock           (clock),           //           clock.clk
		.reset           (reset),           //           reset.reset
		.asmi_busy       (asmi_busy),       //       asmi_busy.asmi_busy
		.asmi_data_valid (asmi_data_valid), // asmi_data_valid.asmi_data_valid
		.asmi_dataout    (asmi_dataout),    //    asmi_dataout.asmi_dataout
		.asmi_addr       (asmi_addr),       //       asmi_addr.asmi_addr
		.asmi_read       (asmi_read),       //       asmi_read.asmi_read
		.asmi_rden       (asmi_rden),       //       asmi_rden.asmi_rden
		.pof_error       (pof_error)        //       pof_error.pof_error
	);

endmodule
